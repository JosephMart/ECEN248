`timescale 1ns / 1ps

module switch_bounce(
    input wire Center,
    output wire J1_0
    );
    
    assign J1_0 = Center;

endmodule
