`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:46:14 11/07/2016 
// Design Name: 
// Module Name:    carry_lookahead_unit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module carry_lookahead_unit(C, G, P, C0);
	 
	 // Ports are wires because we will use dataflow
  output wire [4:1] C; // C4, C3, C2, C1
  input wire [3:0] G, P; // Generates and propagates
  input wire C0; // input carry

  assign #2 C[1] = G[0] | (P[0] & C0);
  assign #2 C[2] = G[1] | (P[1] & G[0]) | (P[1] & P[0] & C0);
  assign #2 C[3] = G[2] | (P[2] & G[1]) | (P[2] & P[1] & G[0]) | (P[2] & P[1] & P[0] & C0);
  assign #2 C[4] = G[3] | (P[3] & G[2]) | (P[3] & P[2] & G[1]) | (P[3] & P[2] & P[1] & G[0]) | (P[3] & P[2] & P[1] & P[0] & C0);
endmodule

//@ladiesmanMB
