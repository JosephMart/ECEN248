`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:13:10 10/24/2016 
// Design Name: 
// Module Name:    adder_2bit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module adder_2bit(Carry, Sum, A, B);
		output wire [1:0] Sum;
		output wire Carry;
		
		input wire [1:0] A;
		input wire [1:0] B;
		wire Cout;
		
		full_adder fa0(Sum[0], Cout, A[0], B[0], 0);
		full_adder fa1(Sum[1], Carry, A[1], B[1], Cout );

endmodule
